class trans;

rand bit ren,wen;
rand logic[15:0] din;
logic [15:0]dout;
bit full, empty;

endclass

